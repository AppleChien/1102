library verilog;
use verilog.vl_types.all;
entity FA_test is
end FA_test;
